interface axi_glb_signal();
    logic clk       ;
    logic rst_n     ;


endinterface