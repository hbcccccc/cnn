module cnn_top_verilog_wrapper2
(
input                                                 clk           ,
input                                                 rst_n         ,
output  wire                                          o_interrupt   ,
output  wire    [23:0]                                o_rgb         ,
output  wire                                          o_rgb_clk     ,
output  wire                                          lcd_de        ,
output  wire                                          lcd_rst_n     ,
output  wire                                          lcd_bl        ,
output  wire                                          lcd_hs        ,
output  wire                                          lcd_vs        ,
output  wire                                          ova_cfg_scl   ,
inout   wire                                          ova_cfg_sda   ,
input   wire                                          i_pclk        ,
input   wire   [7:0]                                  i_data        ,
input   wire                                          href          ,
input   wire                                          vsync         ,

input   [ID_MAX_WIDTH-1           :0]                 arid          ,
input   [ADDR_WIDTH - 1           :0]                 araddr        ,
input   [3                        :0]                 arlen         ,
input   [2                        :0]                 arsize        ,
input   [1                        :0]                 arbrust       ,
input   [1                        :0]                 arlock        ,
input   [3                        :0]                 arcache       ,
input   [2                        :0]                 arprot        ,
input   [3                        :0]                 arqos         ,
input   [3                        :0]                 arregion      ,
input                                                 arvalid       ,
output                                                arready       ,

input   [ID_MAX_WIDTH-1  :0]                          rid           ,
input   [DATA_WIDTH-1    :0]                          rdata         ,
input   [1               :0]                          rresp         ,
input                                                 rlast         ,
input                                                 ruser         ,
input                                                 rvalid        ,
input                                                 rready        ,
input   [ID_MAX_WIDTH-1           :0]                 wid           ,
input   [DATA_WIDTH - 1           :0]                 wdata         ,
input   [DATA_WIDTH/8 -1          :0]                 wstrb         ,
input                                                 wlast         ,
input                                                 wvalid        ,
output                                                wready        ,
input   [ID_MAX_WIDTH-1           :0]                 wid           ,
input   [ADDR_WIDTH - 1           :0]                 waddr         ,
input   [3                        :0]                 wlen          ,
input   [2                        :0]                 wsize         ,
input   [1                        :0]                 wbrust        ,
input   [1                        :0]                 wlock         ,
input   [3                        :0]                 wcache        ,
input   [2                        :0]                 wprot         ,
input   [3                        :0]                 wqos          ,
input                                                 wvalid        ,
output                                                wready        ,
output  [3:0]                                         bid           ,
output  [1:0]                                         bresp         ,
output                                                buser         ,
output                                                bvalid        ,
input                                                 bready     


);

cnn_top_verilog_wrapper inst_cnn_top_verilog_wrapper
(
.clk          (clk              ) ,
.rst_n        (rst_n            ) ,
.o_interrupt  (o_interr         ) ,
.o_rgb        (o_rgb            ) ,
.o_rgb_clk    (o_rgb_cl         ) ,
.lcd_de       (lcd_de           ) ,
.lcd_rst_n    (lcd_rst_n         ) ,
.lcd_bl       (lcd_bl           ) ,
.lcd_hs       (lcd_hs           ) ,
.lcd_vs       (lcd_vs           ) ,
.ova_cfg_scl  (ova_cfg_scl         ) ,
.ova_cfg_sda  (ova_cfg_sda         ) ,
.i_pclk       (i_pclk           ) ,
.i_data       (i_data           ) ,
.href         (href             ) ,
.vsync        (vsync            ) ,
.arid         (arid             ) ,
.araddr       (araddr           ) ,
.arlen        (arlen            ) ,
.arsize       (arsize           ) ,
.arbrust      (arbrust          ) ,
.arlock       (arlock           ) ,
.arcache      (arcache          ) ,
.arprot       (arprot           ) ,
.arqos        (arqos            ) ,
.arregion     (arregion         ) ,
.arvalid      (arvalid          ) ,
.arready      (arready          ) ,
.rid          (rid              ) ,
.rdata        (rdata            ) ,
.rresp        (rresp            ) ,
.rlast        (rlast            ) ,
.ruser        (ruser            ) ,
.rvalid       (rvalid           ) ,
.rready       (rready           ) ,
.wid          (wid              ) ,
.wdata        (wdata            ) ,
.wstrb        (wstrb            ) ,
.wlast        (wlast            ) ,
.wvalid       (wvalid           ) ,
.wready       (wready           ) ,
.wid          (wid              ) ,
.waddr        (waddr            ) ,
.wlen         (wlen             ) ,
.wsize        (wsize            ) ,
.wbrust       (wbrust           ) ,
.wlock        (wlock            ) ,
.wcache       (wcache           ) ,
.wprot        (wprot            ) ,
.wqos         (wqos             ) ,
.wvalid       (wvalid           ) ,
.wready       (wready           ) ,
.bid          (bid              ) ,
.bresp        (bresp            ) ,
.buser        (buser            ) ,
.bvalid       (bvalid           ) ,
.bready       (bready           )
);

endmodule