interface glb_clk_rst          
(
 output bit                  clk   ,    
 output bit                  rst_n
);     

endinterface //intf_sync