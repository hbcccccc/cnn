interface intf_ov7725_data();

logic  pclk;
logic  href;
logic  vsync;
logic [7:0] data;

endinterface