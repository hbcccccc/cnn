interface   intf_i2c;
    wire   sda ;
    wire   scl ;

endinterface